@00000000
13 00 00 00 13 00 00 00 93 00 50 00 13 01 60 00
B3 81 20 00 13 00 00 00 13 00 00 00
