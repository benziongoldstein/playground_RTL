@00000000
13 00 00 00 93 01 00 10 13 01 F0 FF 23 80 21 00
83 80 01 00 03 C2 01 00 13 00 00 00 93 01 40 10
13 01 F0 FF 23 90 21 00 83 90 01 00 03 D2 01 00
13 00 00 00 93 01 80 10 13 01 00 08 23 80 21 00
83 80 01 00 03 C2 01 00 13 00 00 00 93 01 40 10
37 11 00 00 13 01 F1 FF 13 01 11 00 13 01 F1 FF
B7 12 00 00 33 01 51 40 23 90 21 00 83 90 01 00
03 D2 01 00 13 00 00 00 13 00 00 00 73 00 10 00
