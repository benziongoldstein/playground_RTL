@00000000
93 00 50 00 13 01 50 00 93 01 60 00 13 02 40 00
93 02 B0 FF 13 03 A0 FF 93 03 F0 FF 37 04 00 80
63 86 20 00 13 05 10 00 93 05 20 00 13 06 30 00
63 96 30 00 93 06 10 00 13 07 20 00 93 07 30 00
63 46 12 00 13 08 10 00 93 08 20 00 13 09 30 00
63 D6 30 00 93 09 10 00 13 0A 20 00 93 0A 30 00
63 E6 70 00 13 0B 10 00 93 0B 20 00 13 0C 30 00
63 F6 70 00 93 0C 10 00 13 0D 20 00 93 0D 30 00
63 C6 62 00 13 0E 10 00 93 0E 20 00 13 0F 30 00
63 44 54 00 93 0F 10 00 93 02 20 00 13 00 00 00
13 00 00 00 73 00 10 00
