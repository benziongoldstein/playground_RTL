@00000000
13 00 00 00 93 00 60 00 13 01 50 00 B3 81 20 40
13 00 00 00
