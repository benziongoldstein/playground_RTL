@00000000
93 00 50 00 13 01 50 00 93 01 60 00 13 02 40 00
93 02 B0 FF 13 03 A0 FF 93 03 F0 FF 37 04 00 80
63 86 20 00 13 05 10 00 93 05 20 00 13 06 30 00
63 96 30 00 93 06 10 00 13 07 20 00 93 07 30 00
63 46 12 00 13 08 10 00 93 08 20 00 13 09 30 00
13 00 00 00 13 00 00 00 73 00 10 00
