@00000000
13 00 00 00 93 00 50 00 13 01 30 00 B3 E1 20 00
13 02 70 00 93 02 70 00 33 63 52 00 13 00 00 00
