@00000000
13 00 00 00 13 00 00 00 EF 00 80 00 6F 00 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 10 00
23 26 F4 FE 93 07 20 00 23 24 F4 FE 03 27 C4 FE
83 27 84 FE B3 07 F7 00 23 22 F4 FE 03 27 C4 FE
83 27 44 FE B3 07 F7 00 23 20 F4 FE 03 27 84 FE
83 27 04 FE B3 07 F7 00 23 2E F4 FC 03 27 C4 FE
83 27 84 FE B3 07 F7 00 23 22 F4 FE 6F F0 1F FF
